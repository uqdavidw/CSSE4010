    Mac OS X            	   2   �                                           ATTR         �   K                  �     com.apple.lastuseddate#PS       �   ;  com.apple.quarantine ��[    ��    q/0083;5b8c8de8;Slack;77669BAB-220D-42F8-B7E8-70962761C943 